`include "addr_reg_bank_tables.vh"
