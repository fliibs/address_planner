//==========================================================
// Definition of address space TOP_SYS0_IP_A
//==========================================================

`ifndef     ADDR_TOP_SYS0_IP_A
    `define ADDR_TOP_SYS0_IP_A                                       0x0
    `define SIZE_TOP_SYS0_IP_A                                       0x1000
    `define OFFSET_TOP_SYS0_IP_A                                     0x0
`endif

//==========================================================
// Sub address space definition of TOP_SYS0_IP_A
//==========================================================

`ifndef     ADDR_TOP_SYS0_IP_A_MEM_A0
    `define ADDR_TOP_SYS0_IP_A_MEM_A0                                       0x0
    `define SIZE_TOP_SYS0_IP_A_MEM_A0                                       0x400
    `define OFFSET_TOP_SYS0_IP_A_MEM_A0                                     0x0
`endif

`ifndef     ADDR_TOP_SYS0_IP_A_MEM_A1
    `define ADDR_TOP_SYS0_IP_A_MEM_A1                                       0x800
    `define SIZE_TOP_SYS0_IP_A_MEM_A1                                       0x400
    `define OFFSET_TOP_SYS0_IP_A_MEM_A1                                     0x800
`endif
