
//==========================================================
// Definition of reg TOP_SYS0_IP_B_REG_REG0
//==========================================================
#ifndef ADDR_TOP_SYS0_IP_B_REG_REG0
    #define ADDR_TOP_SYS0_IP_B_REG_REG0                                  0x100800
    #define SIZE_TOP_SYS0_IP_B_REG_REG0                                  0x1
    #define OFFSET_TOP_SYS0_IP_B_REG_REG0                                0x0
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD0
    #define OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD0 0
    #define WIDTH_TOP_SYS0_IP_B_REG_REG0_FIELD0  1
    #define MASK_TOP_SYS0_IP_B_REG_REG0_FIELD0   0x1
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD1
    #define OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD1 1
    #define WIDTH_TOP_SYS0_IP_B_REG_REG0_FIELD1  1
    #define MASK_TOP_SYS0_IP_B_REG_REG0_FIELD1   0x2
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD2
    #define OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD2 2
    #define WIDTH_TOP_SYS0_IP_B_REG_REG0_FIELD2  1
    #define MASK_TOP_SYS0_IP_B_REG_REG0_FIELD2   0x4
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD3
    #define OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD3 3
    #define WIDTH_TOP_SYS0_IP_B_REG_REG0_FIELD3  1
    #define MASK_TOP_SYS0_IP_B_REG_REG0_FIELD3   0x8
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD4
    #define OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD4 4
    #define WIDTH_TOP_SYS0_IP_B_REG_REG0_FIELD4  1
    #define MASK_TOP_SYS0_IP_B_REG_REG0_FIELD4   0x10
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD5
    #define OFFSET_TOP_SYS0_IP_B_REG_REG0_FIELD5 5
    #define WIDTH_TOP_SYS0_IP_B_REG_REG0_FIELD5  1
    #define MASK_TOP_SYS0_IP_B_REG_REG0_FIELD5   0x20
#endif


//==========================================================
// Definition of reg TOP_SYS0_IP_B_REG_REG1
//==========================================================
#ifndef ADDR_TOP_SYS0_IP_B_REG_REG1
    #define ADDR_TOP_SYS0_IP_B_REG_REG1                                  0x100801
    #define SIZE_TOP_SYS0_IP_B_REG_REG1                                  0x1
    #define OFFSET_TOP_SYS0_IP_B_REG_REG1                                0x1
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD0
    #define OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD0 0
    #define WIDTH_TOP_SYS0_IP_B_REG_REG1_FIELD0  1
    #define MASK_TOP_SYS0_IP_B_REG_REG1_FIELD0   0x1
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD1
    #define OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD1 1
    #define WIDTH_TOP_SYS0_IP_B_REG_REG1_FIELD1  1
    #define MASK_TOP_SYS0_IP_B_REG_REG1_FIELD1   0x2
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD2
    #define OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD2 2
    #define WIDTH_TOP_SYS0_IP_B_REG_REG1_FIELD2  1
    #define MASK_TOP_SYS0_IP_B_REG_REG1_FIELD2   0x4
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD3
    #define OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD3 3
    #define WIDTH_TOP_SYS0_IP_B_REG_REG1_FIELD3  1
    #define MASK_TOP_SYS0_IP_B_REG_REG1_FIELD3   0x8
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD4
    #define OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD4 4
    #define WIDTH_TOP_SYS0_IP_B_REG_REG1_FIELD4  1
    #define MASK_TOP_SYS0_IP_B_REG_REG1_FIELD4   0x10
#endif

#ifndef OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD5
    #define OFFSET_TOP_SYS0_IP_B_REG_REG1_FIELD5 5
    #define WIDTH_TOP_SYS0_IP_B_REG_REG1_FIELD5  1
    #define MASK_TOP_SYS0_IP_B_REG_REG1_FIELD5   0x20
#endif

